%SYSTEMVAR_DECL
  do_OutHeat1 : BOOL (* Digital Output of Zone x *)
     %DISPLAY_LEVEL 1  %INPUT_LEVEL 16

// Temperature Output 1 Temperature Output Zone 1
;
 do_OutHeat1_stat : BOOL (* status of digital output of Zone x *)
     %INPUT_LEVEL 16

// Status Status Output Zone
;
 do_OutHeat2 : BOOL (* Digital Output of Zone x *)
     %DISPLAY_LEVEL 1  %INPUT_LEVEL 16

// Temperature Output 2 Temperature Output Zone 2
;
 do_OutHeat2_stat : BOOL (* status of digital output of Zone x *)
     %INPUT_LEVEL 16

// Status Status Output Zone
;
 do_OutHeat3 : BOOL (* Digital Output of Zone x *)
     %DISPLAY_LEVEL 1  %INPUT_LEVEL 16

// Temperature Output 3 Temperature Output Zone 3
;
 do_OutHeat3_stat : BOOL (* status of digital output of Zone x *)
     %INPUT_LEVEL 16

// Status Status Output Zone
;
 do_OutHeat4 : BOOL (* Digital Output of Zone x *)
     %DISPLAY_LEVEL 1  %INPUT_LEVEL 16

// Temperature Output 4 Temperature Output Zone 4
;
 do_OutHeat4_stat : BOOL (* status of digital output of Zone x *)
     %INPUT_LEVEL 16

// Status Status Output Zone
;
 do_OutHeat5 : BOOL (* Digital Output of Zone x *)
     %DISPLAY_LEVEL 1  %INPUT_LEVEL 16

// Temperature Output 5 Temperature Output Zone 5
;
 do_OutHeat5_stat : BOOL (* status of digital output of Zone x *)
     %INPUT_LEVEL 16

// Status Status Output Zone
;
 do_OutHeat6 : BOOL (* Digital Output of Zone x *)
     %DISPLAY_LEVEL 1  %INPUT_LEVEL 16

// Temperature Output 6 Temperature Output Zone 6
;
 do_OutHeat6_stat : BOOL (* status of digital output of Zone x *)
     %INPUT_LEVEL 16

// Status Status Output Zone
;
 do_OutHeat7 : BOOL (* Digital Output of Zone x *)
     %DISPLAY_LEVEL 1  %INPUT_LEVEL 16

// Temperature Output 7 Temperature Output Zone 7
;
 do_OutHeat7_stat : BOOL (* status of digital output of Zone x *)
     %INPUT_LEVEL 16

// Status Status Output Zone
;
 do_OutHeat8 : BOOL (* Digital Output of Zone x *)
     %DISPLAY_LEVEL 1  %INPUT_LEVEL 16

// Temperature Output 8 Temperature Output Zone 8
;
 do_OutHeat8_stat : BOOL (* status of digital output of Zone x *)
     %INPUT_LEVEL 16

// Status Status Output Zone
;
 do_OutHeat9 : BOOL (* Digital Output of Zone x *)
     %DISPLAY_LEVEL 1  %INPUT_LEVEL 16

// Temperature Output 9 Temperature Output Zone 9
;
 do_OutHeat9_stat : BOOL (* status of digital output of Zone x *)
     %INPUT_LEVEL 16

// Status Status Output Zone
;
 do_OutHeat10 : BOOL (* Digital Output of Zone x *)
     %DISPLAY_LEVEL 1  %INPUT_LEVEL 16

// Temperature Output 10 Temperature Output Zone 10
;
 do_OutHeat10_stat : BOOL (* status of digital output of Zone x *)
     %INPUT_LEVEL 16

// Status Status Output Zone
;
 do_OutHeat11 : BOOL (* Digital Output of Zone x *)
     %DISPLAY_LEVEL 1  %INPUT_LEVEL 16

// Temperature Output 11 Temperature Output Zone 11
;
 do_OutHeat11_stat : BOOL (* status of digital output of Zone x *)
     %INPUT_LEVEL 16

// Status Status Output Zone
;
 do_OutHeat12 : BOOL (* Digital Output of Zone x *)
     %DISPLAY_LEVEL 1  %INPUT_LEVEL 16

// Temperature Output 12 Temperature Output Zone 12
;
 do_OutHeat12_stat : BOOL (* status of digital output of Zone x *)
     %INPUT_LEVEL 16

// Status Status Output Zone
;
%END



#END_OF_IEC_PART

@Puma @IecEditor 6 60 @Sve 25 
@@@BEG_Comment@@@

@@@END_Comment@@@

@BEG_Contents 

@BEG_Export 
@RT(16)SveTreeContainer 
24 
@SysVar @RT(11)do_OutHeat1 @RT(0) @T @F @DT @RT(4)BOOL @RT(0) @T @T @BASIC 0 @F 
@F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(24)Digital Output of Zone x 
@RT(1)1 @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(20)Temperature Output 1 @RT(25)Temperature Output Zone 1 @RT(0) @RT(0) @RT(0) 
@END_Attrib 
1 
@AttrSym @RT(11)do_OutHeat1 @RT(0) @F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(24)Digital Output of Zone x 
@RT(1)1 @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(20)Temperature Output 1 @RT(25)Temperature Output Zone 1 @RT(0) @RT(0) @RT(0) 
@END_Attrib 


@SysVar @RT(16)do_OutHeat1_stat @RT(0) @T @F @DT @RT(4)BOOL @RT(0) @T @T @BASIC 0 @F 
@F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(34)status of digital output of Zone x 
@RT(0) @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(6)Status @RT(18)Status Output Zone @RT(0) @RT(0) @RT(0) 
@END_Attrib 
1 
@AttrSym @RT(16)do_OutHeat1_stat @RT(0) @F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(34)status of digital output of Zone x 
@RT(0) @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(6)Status @RT(18)Status Output Zone @RT(0) @RT(0) @RT(0) 
@END_Attrib 


@SysVar @RT(11)do_OutHeat2 @RT(0) @T @F @DT @RT(4)BOOL @RT(0) @T @T @BASIC 0 @F 
@F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(24)Digital Output of Zone x 
@RT(1)1 @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(20)Temperature Output 2 @RT(25)Temperature Output Zone 2 @RT(0) @RT(0) @RT(0) 
@END_Attrib 
1 
@AttrSym @RT(11)do_OutHeat2 @RT(0) @F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(24)Digital Output of Zone x 
@RT(1)1 @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(20)Temperature Output 2 @RT(25)Temperature Output Zone 2 @RT(0) @RT(0) @RT(0) 
@END_Attrib 


@SysVar @RT(16)do_OutHeat2_stat @RT(0) @T @F @DT @RT(4)BOOL @RT(0) @T @T @BASIC 0 @F 
@F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(34)status of digital output of Zone x 
@RT(0) @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(6)Status @RT(18)Status Output Zone @RT(0) @RT(0) @RT(0) 
@END_Attrib 
1 
@AttrSym @RT(16)do_OutHeat2_stat @RT(0) @F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(34)status of digital output of Zone x 
@RT(0) @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(6)Status @RT(18)Status Output Zone @RT(0) @RT(0) @RT(0) 
@END_Attrib 


@SysVar @RT(11)do_OutHeat3 @RT(0) @T @F @DT @RT(4)BOOL @RT(0) @T @T @BASIC 0 @F 
@F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(24)Digital Output of Zone x 
@RT(1)1 @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(20)Temperature Output 3 @RT(25)Temperature Output Zone 3 @RT(0) @RT(0) @RT(0) 
@END_Attrib 
1 
@AttrSym @RT(11)do_OutHeat3 @RT(0) @F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(24)Digital Output of Zone x 
@RT(1)1 @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(20)Temperature Output 3 @RT(25)Temperature Output Zone 3 @RT(0) @RT(0) @RT(0) 
@END_Attrib 


@SysVar @RT(16)do_OutHeat3_stat @RT(0) @T @F @DT @RT(4)BOOL @RT(0) @T @T @BASIC 0 @F 
@F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(34)status of digital output of Zone x 
@RT(0) @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(6)Status @RT(18)Status Output Zone @RT(0) @RT(0) @RT(0) 
@END_Attrib 
1 
@AttrSym @RT(16)do_OutHeat3_stat @RT(0) @F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(34)status of digital output of Zone x 
@RT(0) @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(6)Status @RT(18)Status Output Zone @RT(0) @RT(0) @RT(0) 
@END_Attrib 


@SysVar @RT(11)do_OutHeat4 @RT(0) @T @F @DT @RT(4)BOOL @RT(0) @T @T @BASIC 0 @F 
@F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(24)Digital Output of Zone x 
@RT(1)1 @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(20)Temperature Output 4 @RT(25)Temperature Output Zone 4 @RT(0) @RT(0) @RT(0) 
@END_Attrib 
1 
@AttrSym @RT(11)do_OutHeat4 @RT(0) @F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(24)Digital Output of Zone x 
@RT(1)1 @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(20)Temperature Output 4 @RT(25)Temperature Output Zone 4 @RT(0) @RT(0) @RT(0) 
@END_Attrib 


@SysVar @RT(16)do_OutHeat4_stat @RT(0) @T @F @DT @RT(4)BOOL @RT(0) @T @T @BASIC 0 @F 
@F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(34)status of digital output of Zone x 
@RT(0) @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(6)Status @RT(18)Status Output Zone @RT(0) @RT(0) @RT(0) 
@END_Attrib 
1 
@AttrSym @RT(16)do_OutHeat4_stat @RT(0) @F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(34)status of digital output of Zone x 
@RT(0) @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(6)Status @RT(18)Status Output Zone @RT(0) @RT(0) @RT(0) 
@END_Attrib 


@SysVar @RT(11)do_OutHeat5 @RT(0) @T @F @DT @RT(4)BOOL @RT(0) @T @T @BASIC 0 @F 
@F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(24)Digital Output of Zone x 
@RT(1)1 @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(20)Temperature Output 5 @RT(25)Temperature Output Zone 5 @RT(0) @RT(0) @RT(0) 
@END_Attrib 
1 
@AttrSym @RT(11)do_OutHeat5 @RT(0) @F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(24)Digital Output of Zone x 
@RT(1)1 @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(20)Temperature Output 5 @RT(25)Temperature Output Zone 5 @RT(0) @RT(0) @RT(0) 
@END_Attrib 


@SysVar @RT(16)do_OutHeat5_stat @RT(0) @T @F @DT @RT(4)BOOL @RT(0) @T @T @BASIC 0 @F 
@F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(34)status of digital output of Zone x 
@RT(0) @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(6)Status @RT(18)Status Output Zone @RT(0) @RT(0) @RT(0) 
@END_Attrib 
1 
@AttrSym @RT(16)do_OutHeat5_stat @RT(0) @F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(34)status of digital output of Zone x 
@RT(0) @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(6)Status @RT(18)Status Output Zone @RT(0) @RT(0) @RT(0) 
@END_Attrib 


@SysVar @RT(11)do_OutHeat6 @RT(0) @T @F @DT @RT(4)BOOL @RT(0) @T @T @BASIC 0 @F 
@F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(24)Digital Output of Zone x 
@RT(1)1 @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(20)Temperature Output 6 @RT(25)Temperature Output Zone 6 @RT(0) @RT(0) @RT(0) 
@END_Attrib 
1 
@AttrSym @RT(11)do_OutHeat6 @RT(0) @F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(24)Digital Output of Zone x 
@RT(1)1 @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(20)Temperature Output 6 @RT(25)Temperature Output Zone 6 @RT(0) @RT(0) @RT(0) 
@END_Attrib 


@SysVar @RT(16)do_OutHeat6_stat @RT(0) @T @F @DT @RT(4)BOOL @RT(0) @T @T @BASIC 0 @F 
@F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(34)status of digital output of Zone x 
@RT(0) @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(6)Status @RT(18)Status Output Zone @RT(0) @RT(0) @RT(0) 
@END_Attrib 
1 
@AttrSym @RT(16)do_OutHeat6_stat @RT(0) @F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(34)status of digital output of Zone x 
@RT(0) @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(6)Status @RT(18)Status Output Zone @RT(0) @RT(0) @RT(0) 
@END_Attrib 


@SysVar @RT(11)do_OutHeat7 @RT(0) @T @F @DT @RT(4)BOOL @RT(0) @T @T @BASIC 0 @F 
@F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(24)Digital Output of Zone x 
@RT(1)1 @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(20)Temperature Output 7 @RT(25)Temperature Output Zone 7 @RT(0) @RT(0) @RT(0) 
@END_Attrib 
1 
@AttrSym @RT(11)do_OutHeat7 @RT(0) @F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(24)Digital Output of Zone x 
@RT(1)1 @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(20)Temperature Output 7 @RT(25)Temperature Output Zone 7 @RT(0) @RT(0) @RT(0) 
@END_Attrib 


@SysVar @RT(16)do_OutHeat7_stat @RT(0) @T @F @DT @RT(4)BOOL @RT(0) @T @T @BASIC 0 @F 
@F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(34)status of digital output of Zone x 
@RT(0) @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(6)Status @RT(18)Status Output Zone @RT(0) @RT(0) @RT(0) 
@END_Attrib 
1 
@AttrSym @RT(16)do_OutHeat7_stat @RT(0) @F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(34)status of digital output of Zone x 
@RT(0) @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(6)Status @RT(18)Status Output Zone @RT(0) @RT(0) @RT(0) 
@END_Attrib 


@SysVar @RT(11)do_OutHeat8 @RT(0) @T @F @DT @RT(4)BOOL @RT(0) @T @T @BASIC 0 @F 
@F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(24)Digital Output of Zone x 
@RT(1)1 @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(20)Temperature Output 8 @RT(25)Temperature Output Zone 8 @RT(0) @RT(0) @RT(0) 
@END_Attrib 
1 
@AttrSym @RT(11)do_OutHeat8 @RT(0) @F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(24)Digital Output of Zone x 
@RT(1)1 @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(20)Temperature Output 8 @RT(25)Temperature Output Zone 8 @RT(0) @RT(0) @RT(0) 
@END_Attrib 


@SysVar @RT(16)do_OutHeat8_stat @RT(0) @T @F @DT @RT(4)BOOL @RT(0) @T @T @BASIC 0 @F 
@F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(34)status of digital output of Zone x 
@RT(0) @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(6)Status @RT(18)Status Output Zone @RT(0) @RT(0) @RT(0) 
@END_Attrib 
1 
@AttrSym @RT(16)do_OutHeat8_stat @RT(0) @F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(34)status of digital output of Zone x 
@RT(0) @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(6)Status @RT(18)Status Output Zone @RT(0) @RT(0) @RT(0) 
@END_Attrib 


@SysVar @RT(11)do_OutHeat9 @RT(0) @T @F @DT @RT(4)BOOL @RT(0) @T @T @BASIC 0 @F 
@F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(24)Digital Output of Zone x 
@RT(1)1 @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(20)Temperature Output 9 @RT(25)Temperature Output Zone 9 @RT(0) @RT(0) @RT(0) 
@END_Attrib 
1 
@AttrSym @RT(11)do_OutHeat9 @RT(0) @F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(24)Digital Output of Zone x 
@RT(1)1 @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(20)Temperature Output 9 @RT(25)Temperature Output Zone 9 @RT(0) @RT(0) @RT(0) 
@END_Attrib 


@SysVar @RT(16)do_OutHeat9_stat @RT(0) @T @F @DT @RT(4)BOOL @RT(0) @T @T @BASIC 0 @F 
@F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(34)status of digital output of Zone x 
@RT(0) @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(6)Status @RT(18)Status Output Zone @RT(0) @RT(0) @RT(0) 
@END_Attrib 
1 
@AttrSym @RT(16)do_OutHeat9_stat @RT(0) @F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(34)status of digital output of Zone x 
@RT(0) @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(6)Status @RT(18)Status Output Zone @RT(0) @RT(0) @RT(0) 
@END_Attrib 


@SysVar @RT(12)do_OutHeat10 @RT(0) @T @F @DT @RT(4)BOOL @RT(0) @T @T @BASIC 0 @F 
@F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(24)Digital Output of Zone x 
@RT(1)1 @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(21)Temperature Output 10 @RT(26)Temperature Output Zone 10 @RT(0) @RT(0) @RT(0) 
@END_Attrib 
1 
@AttrSym @RT(12)do_OutHeat10 @RT(0) @F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(24)Digital Output of Zone x 
@RT(1)1 @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(21)Temperature Output 10 @RT(26)Temperature Output Zone 10 @RT(0) @RT(0) @RT(0) 
@END_Attrib 


@SysVar @RT(17)do_OutHeat10_stat @RT(0) @T @F @DT @RT(4)BOOL @RT(0) @T @T @BASIC 0 @F 
@F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(34)status of digital output of Zone x 
@RT(0) @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(6)Status @RT(18)Status Output Zone @RT(0) @RT(0) @RT(0) 
@END_Attrib 
1 
@AttrSym @RT(17)do_OutHeat10_stat @RT(0) @F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(34)status of digital output of Zone x 
@RT(0) @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(6)Status @RT(18)Status Output Zone @RT(0) @RT(0) @RT(0) 
@END_Attrib 


@SysVar @RT(12)do_OutHeat11 @RT(0) @T @F @DT @RT(4)BOOL @RT(0) @T @T @BASIC 0 @F 
@F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(24)Digital Output of Zone x 
@RT(1)1 @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(21)Temperature Output 11 @RT(26)Temperature Output Zone 11 @RT(0) @RT(0) @RT(0) 
@END_Attrib 
1 
@AttrSym @RT(12)do_OutHeat11 @RT(0) @F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(24)Digital Output of Zone x 
@RT(1)1 @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(21)Temperature Output 11 @RT(26)Temperature Output Zone 11 @RT(0) @RT(0) @RT(0) 
@END_Attrib 


@SysVar @RT(17)do_OutHeat11_stat @RT(0) @T @F @DT @RT(4)BOOL @RT(0) @T @T @BASIC 0 @F 
@F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(34)status of digital output of Zone x 
@RT(0) @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(6)Status @RT(18)Status Output Zone @RT(0) @RT(0) @RT(0) 
@END_Attrib 
1 
@AttrSym @RT(17)do_OutHeat11_stat @RT(0) @F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(34)status of digital output of Zone x 
@RT(0) @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(6)Status @RT(18)Status Output Zone @RT(0) @RT(0) @RT(0) 
@END_Attrib 


@SysVar @RT(12)do_OutHeat12 @RT(0) @T @F @DT @RT(4)BOOL @RT(0) @T @T @BASIC 0 @F 
@F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(24)Digital Output of Zone x 
@RT(1)1 @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(21)Temperature Output 12 @RT(26)Temperature Output Zone 12 @RT(0) @RT(0) @RT(0) 
@END_Attrib 
1 
@AttrSym @RT(12)do_OutHeat12 @RT(0) @F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(24)Digital Output of Zone x 
@RT(1)1 @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(21)Temperature Output 12 @RT(26)Temperature Output Zone 12 @RT(0) @RT(0) @RT(0) 
@END_Attrib 


@SysVar @RT(17)do_OutHeat12_stat @RT(0) @T @F @DT @RT(4)BOOL @RT(0) @T @T @BASIC 0 @F 
@F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(34)status of digital output of Zone x 
@RT(0) @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(6)Status @RT(18)Status Output Zone @RT(0) @RT(0) @RT(0) 
@END_Attrib 
1 
@AttrSym @RT(17)do_OutHeat12_stat @RT(0) @F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(34)status of digital output of Zone x 
@RT(0) @RT(2)16 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(6)Status @RT(18)Status Output Zone @RT(0) @RT(0) @RT(0) 
@END_Attrib 


@RT(15)SETreeContainer 
0 
@RT(15)SOTreeContainer 
0 

@RT(15)SATreeContainer 
0 

@RT(21)SExtAttrTreeContainer 
0 
@END_Export 

@END_Contents 
