%SYSTEMVAR_DECL
  di_EmergencyStop1 : BOOL
     %DISPLAY_LEVEL 1 
// DI Emergency stop 1 DI emergency stop 1
;
 di_EmergencyStop1_stat : BOOL
    
// Emergency stop 1 state DI emergency stop 1 state
;
 di_EmergencyStop2 : BOOL
     %DISPLAY_LEVEL 1 
// DI Emergency stop 2 DI emergency stop 2
;
 di_EmergencyStop2_stat : BOOL
    
// Emergency stop 2 state DI emergency stop 2 state
;
 di_EmergencyStop3 : BOOL
     %DISPLAY_LEVEL 1 
// DI Emergency stop 3 DI emergency stop 3
;
 di_EmergencyStop3_stat : BOOL
    
// Emergency stop 3 state DI emergency stop 3 state
;
 di_EmergencyStop4 : BOOL
     %DISPLAY_LEVEL 1 
// DI Emergency stop 4 DI emergency stop 4
;
 di_EmergencyStop4_stat : BOOL
    
// Emergency stop 4 state DI emergency stop 4 state
;
%END



#END_OF_IEC_PART

@Puma @IecEditor 6 97 @Sve 25 
@@@BEG_Comment@@@

@@@END_Comment@@@

@BEG_Contents 

@BEG_Export 
@RT(16)SveTreeContainer 
8 
@SysVar @RT(17)di_EmergencyStop1 @RT(0) @T @F @DT @RT(4)BOOL @RT(0) @T @T @BASIC 0 @F 
@F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(0) 
@RT(1)1 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(19)DI Emergency stop 1 @RT(19)DI emergency stop 1 @RT(0) @RT(0) @RT(0) 
@END_Attrib 
1 
@AttrSym @RT(17)di_EmergencyStop1 @RT(0) @F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(0) 
@RT(1)1 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(19)DI Emergency stop 1 @RT(19)DI emergency stop 1 @RT(0) @RT(0) @RT(0) 
@END_Attrib 


@SysVar @RT(22)di_EmergencyStop1_stat @RT(0) @T @F @DT @RT(4)BOOL @RT(0) @T @T @BASIC 0 @F 
@F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(22)Emergency stop 1 state @RT(25)DI emergency stop 1 state @RT(0) @RT(0) @RT(0) 
@END_Attrib 
1 
@AttrSym @RT(22)di_EmergencyStop1_stat @RT(0) @F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(22)Emergency stop 1 state @RT(25)DI emergency stop 1 state @RT(0) @RT(0) @RT(0) 
@END_Attrib 


@SysVar @RT(17)di_EmergencyStop2 @RT(0) @T @F @DT @RT(4)BOOL @RT(0) @T @T @BASIC 0 @F 
@F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(0) 
@RT(1)1 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(19)DI Emergency stop 2 @RT(19)DI emergency stop 2 @RT(0) @RT(0) @RT(0) 
@END_Attrib 
1 
@AttrSym @RT(17)di_EmergencyStop2 @RT(0) @F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(0) 
@RT(1)1 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(19)DI Emergency stop 2 @RT(19)DI emergency stop 2 @RT(0) @RT(0) @RT(0) 
@END_Attrib 


@SysVar @RT(22)di_EmergencyStop2_stat @RT(0) @T @F @DT @RT(4)BOOL @RT(0) @T @T @BASIC 0 @F 
@F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(22)Emergency stop 2 state @RT(25)DI emergency stop 2 state @RT(0) @RT(0) @RT(0) 
@END_Attrib 
1 
@AttrSym @RT(22)di_EmergencyStop2_stat @RT(0) @F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(22)Emergency stop 2 state @RT(25)DI emergency stop 2 state @RT(0) @RT(0) @RT(0) 
@END_Attrib 


@SysVar @RT(17)di_EmergencyStop3 @RT(0) @T @F @DT @RT(4)BOOL @RT(0) @T @T @BASIC 0 @F 
@F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(0) 
@RT(1)1 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(19)DI Emergency stop 3 @RT(19)DI emergency stop 3 @RT(0) @RT(0) @RT(0) 
@END_Attrib 
1 
@AttrSym @RT(17)di_EmergencyStop3 @RT(0) @F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(0) 
@RT(1)1 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(19)DI Emergency stop 3 @RT(19)DI emergency stop 3 @RT(0) @RT(0) @RT(0) 
@END_Attrib 


@SysVar @RT(22)di_EmergencyStop3_stat @RT(0) @T @F @DT @RT(4)BOOL @RT(0) @T @T @BASIC 0 @F 
@F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(22)Emergency stop 3 state @RT(25)DI emergency stop 3 state @RT(0) @RT(0) @RT(0) 
@END_Attrib 
1 
@AttrSym @RT(22)di_EmergencyStop3_stat @RT(0) @F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(22)Emergency stop 3 state @RT(25)DI emergency stop 3 state @RT(0) @RT(0) @RT(0) 
@END_Attrib 


@SysVar @RT(17)di_EmergencyStop4 @RT(0) @T @F @DT @RT(4)BOOL @RT(0) @T @T @BASIC 0 @F 
@F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(0) 
@RT(1)1 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(19)DI Emergency stop 4 @RT(19)DI emergency stop 4 @RT(0) @RT(0) @RT(0) 
@END_Attrib 
1 
@AttrSym @RT(17)di_EmergencyStop4 @RT(0) @F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(0) 
@RT(1)1 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(19)DI Emergency stop 4 @RT(19)DI emergency stop 4 @RT(0) @RT(0) @RT(0) 
@END_Attrib 


@SysVar @RT(22)di_EmergencyStop4_stat @RT(0) @T @F @DT @RT(4)BOOL @RT(0) @T @T @BASIC 0 @F 
@F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(22)Emergency stop 4 state @RT(25)DI emergency stop 4 state @RT(0) @RT(0) @RT(0) 
@END_Attrib 
1 
@AttrSym @RT(22)di_EmergencyStop4_stat @RT(0) @F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(22)Emergency stop 4 state @RT(25)DI emergency stop 4 state @RT(0) @RT(0) @RT(0) 
@END_Attrib 


@RT(15)SETreeContainer 
0 
@RT(15)SOTreeContainer 
0 

@RT(15)SATreeContainer 
0 

@RT(21)SExtAttrTreeContainer 
0 
@END_Export 

@END_Contents 
