%SYSTEMVAR_DECL
  di_Open : BOOL
     %DISPLAY_LEVEL 1 
// DI sg mold open DI safety gate mold open
;
 di_Open_stat : BOOL
    
// DI open state DI safety gate open
;
 di_Closed : BOOL
     %DISPLAY_LEVEL 1 
// DI sg mold closed DI safety gate mold closed
;
 di_Closed_stat : BOOL
    
// DI closed state DI safety gate closed state
;
%END



#END_OF_IEC_PART

@Puma @IecEditor 6 97 @Sve 25 
@@@BEG_Comment@@@

@@@END_Comment@@@

@BEG_Contents 

@BEG_Export 
@RT(16)SveTreeContainer 
4 
@SysVar @RT(7)di_Open @RT(0) @T @F @DT @RT(4)BOOL @RT(0) @T @T @BASIC 0 @F 
@F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(0) 
@RT(1)1 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(15)DI sg mold open @RT(24)DI safety gate mold open @RT(0) @RT(0) @RT(0) 
@END_Attrib 
1 
@AttrSym @RT(7)di_Open @RT(0) @F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(0) 
@RT(1)1 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(15)DI sg mold open @RT(24)DI safety gate mold open @RT(0) @RT(0) @RT(0) 
@END_Attrib 


@SysVar @RT(12)di_Open_stat @RT(0) @T @F @DT @RT(4)BOOL @RT(0) @T @T @BASIC 0 @F 
@F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(13)DI open state @RT(19)DI safety gate open @RT(0) @RT(0) @RT(0) 
@END_Attrib 
1 
@AttrSym @RT(12)di_Open_stat @RT(0) @F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(13)DI open state @RT(19)DI safety gate open @RT(0) @RT(0) @RT(0) 
@END_Attrib 


@SysVar @RT(9)di_Closed @RT(0) @T @F @DT @RT(4)BOOL @RT(0) @T @T @BASIC 0 @F 
@F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(0) 
@RT(1)1 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(17)DI sg mold closed @RT(26)DI safety gate mold closed @RT(0) @RT(0) @RT(0) 
@END_Attrib 
1 
@AttrSym @RT(9)di_Closed @RT(0) @F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(0) 
@RT(1)1 @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(17)DI sg mold closed @RT(26)DI safety gate mold closed @RT(0) @RT(0) @RT(0) 
@END_Attrib 


@SysVar @RT(14)di_Closed_stat @RT(0) @T @F @DT @RT(4)BOOL @RT(0) @T @T @BASIC 0 @F 
@F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(15)DI closed state @RT(27)DI safety gate closed state @RT(0) @RT(0) @RT(0) 
@END_Attrib 
1 
@AttrSym @RT(14)di_Closed_stat @RT(0) @F @F 
@T 
@BEG_Attrib 
4 @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) @RT(0) 
@RT(15)DI closed state @RT(27)DI safety gate closed state @RT(0) @RT(0) @RT(0) 
@END_Attrib 


@RT(15)SETreeContainer 
0 
@RT(15)SOTreeContainer 
0 

@RT(15)SATreeContainer 
0 

@RT(21)SExtAttrTreeContainer 
0 
@END_Export 

@END_Contents 
