%IMPORT_OVER_LISTFILE_OBJECT
 tevUpdateEventNotification
, tevRequestEventNotification

END_IMPORT

%SYSTEMEVENT_DECL
  evUpdateEventNotification : tevUpdateEventNotification
;
 evRequestEventNotification : tevRequestEventNotification
;
%END



#END_OF_IEC_PART

@Puma @IecEditor 6 131 @Sve 25 
@@@BEG_Comment@@@

@@@END_Comment@@@

@BEG_Contents 

@BEG_Export 
@RT(16)SveTreeContainer 
0 
@RT(15)SETreeContainer 
2 
@SysEvent @RT(25)evUpdateEventNotification @RT(0) @T @T @DERIVED 0 @F @RT(26)tevUpdateEventNotification @F 
@T 
@BEG_Attrib 
13 @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) 
@END_Attrib 
0 


@SysEvent @RT(26)evRequestEventNotification @RT(0) @T @T @DERIVED 0 @F @RT(27)tevRequestEventNotification @F 
@T 
@BEG_Attrib 
13 @RT(0) @RT(0) 
@RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) @RT(0) 
@RT(0) 
@END_Attrib 
0 


@RT(15)SOTreeContainer 
0 

@RT(15)SATreeContainer 
0 

@RT(21)SExtAttrTreeContainer 
0 
@END_Export 

@END_Contents 
