%SYSTEM_ALARM
  erRetainVarSupervision
 %CLASS 3 %ACKNOWLEDGEMENT %USER_AND_APPLICATION %PROTOCOL %YES

// Writing retain-variables exceeded limit!
 ;
%END



#END_OF_IEC_PART

@Puma @IecEditor 6 159 @Sve 25 
@@@BEG_Comment@@@

@@@END_Comment@@@

@BEG_Contents 

@BEG_Export 
@RT(16)SveTreeContainer 
0 
@RT(15)SETreeContainer 
0 
@RT(15)SOTreeContainer 
0 

@RT(15)SATreeContainer 
1 @BEG_Attrib 
15 @RT(0) @RT(0) 
@RT(22)erRetainVarSupervision @RT(1)3 @RT(1)y @RT(0) @RT(0) @RT(20)User and Application @RT(40)Writing retain-variables exceeded limit! 
@END_Attrib 
@F 


@RT(21)SExtAttrTreeContainer 
0 
@END_Export 

@END_Contents 
